`include "/MDSD/Extra_credit_sessions/Verilogreview/DisplayComp.v";

module testbench;
    reg [3:0] A=0, B=0;
    reg clk=0;
    wire [6:0] SegmentData;
    top UUT


    endmodule